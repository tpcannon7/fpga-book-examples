module binary_decoder (
    input logic [ 3:0] in,
    input logic [15:0] out
);


endmodule
